module wrapper_MISR #( 
	parameter int unsigned NBIT_DATA = 64,
	parameter int unsigned NBIT_ADDR = 64,
	parameter int unsigned NBIT_REGS = 64, 
	parameter int unsigned START_ADDR = 2**25
	)(
	input 	logic 					clk_i,   
	input 	logic 					rst_ni, 
	input	logic 					req_i,
	input	logic					we_i,
	input 	logic [NBIT_DATA-1:0]	data_i,
	input 	logic [NBIT_ADDR-1:0]	addr_i,
	output 	logic [NBIT_DATA-1:0]	data_o	
);

	//ADDRESSES OF THE CONTROL REGISTERS
	localparam MISR_PERIPH_START_ADDR 				= START_ADDR; //64'h0000000002000000 --> from 2^25, which is the size of the SRAM
	localparam MISR_CONTROL_CONTROL_REG_OFFSET 		= 64'h0000000000000000;
	localparam MISR_CONTROL_COEFFICIENTS_REG_OFFSET	= 64'h0000000000000040;
	localparam MISR_CONTROL_SIGNATURE_REG_OFFSET 	= 64'h0000000000000080;
	localparam MISR_CONTROL_DONE_REG_OFFSET			= 64'h00000000000000C0;

	localparam int MISR_CONTROL_ENABLE_BIT 			= 0;
	localparam int MISR_CONTROL_RESET_BIT 			= 1;
	localparam int MISR_CONTROL_DONE_IN_BIT 		= 2;

	localparam MISR_CONTROL_CONTROL_REG_ADDR 		= MISR_PERIPH_START_ADDR + MISR_CONTROL_CONTROL_REG_OFFSET;
	localparam MISR_CONTROL_COEFFICIENTS_REG_ADDR	= MISR_PERIPH_START_ADDR + MISR_CONTROL_COEFFICIENTS_REG_OFFSET;
	localparam MISR_CONTROL_SIGNATURE_REG_ADDR		= MISR_PERIPH_START_ADDR + MISR_CONTROL_SIGNATURE_REG_OFFSET;
	localparam MISR_CONTROL_DONE_REG_ADDR			= MISR_PERIPH_START_ADDR + MISR_CONTROL_DONE_REG_OFFSET;

	logic en_MISR, rst_MISR;
	logic done_bit;
	logic [NBIT_REGS-1:0] control_reg_in, control_reg_out;
	logic [NBIT_REGS-1:0] coeff_reg_in, coeff_reg_out;
	logic [NBIT_REGS-1:0] signature_reg_in, signature_reg_out;
	logic [NBIT_REGS-1:0] done_reg_in, done_reg_out;

	
	// control register, contains enable and reset bits    
	// SW: rw permission
	// HW: ro permission
	control_reg  #(
		.NBIT(NBIT_REGS)
	) control_register (
		.clk(clk_i), .rst_n(rst_ni), .d(control_reg_in), .q(control_reg_out)
	);
	// coefficients register   
	// SW: rw permission
	// HW: ro permission  
	control_reg  #(
		.NBIT(NBIT_REGS)
	) coefficient_register (
		.clk(clk_i), .rst_n(rst_ni), .d(coeff_reg_in), .q(coeff_reg_out)
	);
	// signature register
	// SW: ro permission
	// HW: rw permission
	control_reg  #(
		.NBIT(NBIT_REGS)
	) signature_register (
		.clk(clk_i), .rst_n(rst_ni), .d(signature_reg_in), .q(signature_reg_out)
	);
	// done bit register (32bits register due to byte alignment)
	// SW: ro permission
	// HW: rw permission
	control_reg  #(
		.NBIT(NBIT_REGS)
	) done_register (
		.clk(clk_i), .rst_n(rst_MISR), .d(done_reg_in), .q(done_reg_out)
	); 

	//MISR
	generic_MISR #(
		.N (NBIT_DATA)
	) MISR (
		.clk 		(clk_i),
		.rst_n 		(rst_MISR),
		.datain 	(data_i),
		.en 		(en_MISR),
		.done_in 	(control_reg_out[MISR_CONTROL_DONE_IN_BIT]),
		.coeff 		(coeff_reg_out),
		.out_sig 	(signature_reg_in), //output
		.done_out 	(done_bit) //output
	);

	always_comb begin 
		//initialize all register input signals
		rst_MISR = rst_ni | control_reg_in[MISR_CONTROL_RESET_BIT];
		en_MISR = control_reg_in[MISR_CONTROL_ENABLE_BIT];
		control_reg_in = control_reg_out;
		coeff_reg_in = coeff_reg_out;
		done_reg_in = {{(NBIT_REGS-1){1'b0}} , done_bit};
		data_o = '0; //if a read request is not specified, simply put all 0 in output (it will be ignored by the bus anyway)

		if (req_i == 1'b1) begin
			// check if the transaction on the AXI bus is towards the MISR registers
			case (addr_i)
				//control register
				MISR_CONTROL_CONTROL_REG_ADDR : begin 
					if (we_i == 1'b1) begin
						control_reg_in = data_i;
					end
					else begin
						data_o = control_reg_out;
					end
				end
				//coefficients register
				MISR_CONTROL_COEFFICIENTS_REG_ADDR : begin
					if (we_i == 1'b1) begin
						coeff_reg_in = data_i;
					end
					else begin
						data_o = coeff_reg_out;
					end
				end
				//signature register
				MISR_CONTROL_SIGNATURE_REG_ADDR : begin
					//this register can only be written by the MISR
					//so, if a write request is issued, nothing will happen
					if (we_i == 1'b0) begin
						data_o = signature_reg_out;
					end
				end
				//done register
				MISR_CONTROL_DONE_REG_ADDR : begin
					//this register can only be written by the MISR
					//so, if a write request is issued, nothing will happen
					if (we_i == 1'b0) begin
						data_o = done_reg_out;
					end
				end
				default : data_o = '0;
			endcase
		end
		
		
	end

endmodule : wrapper_MISR
